LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.numeric_std.ALL;

ENTITY WR_BLOCK IS
	PORT (
		clk : IN STD_LOGIC;
		rst : IN STD_LOGIC;
		ready_w : OUT STD_LOGIC;
		valid_r : IN STD_LOGIC;
		data_in : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		sub_data_in : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		load_adr_in : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		-- memory
		adres_memory : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        memory_data : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        question_memory : OUT STD_LOGIC;
        memory_data_ready : IN STD_LOGIC;
		-- registers
		adres_registers : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        registers_data : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        question_registers : OUT STD_LOGIC;
        registers_data_ready : IN STD_LOGIC
	);
END WR_BLOCK;

ARCHITECTURE rtl OF WR_BLOCK IS

BEGIN
	main : PROCESS (clk, rst)

		VARIABLE valid_map : STD_LOGIC;
		VARIABLE ready_map : STD_LOGIC;
		VARIABLE data : STD_LOGIC_VECTOR(3 DOWNTO 0);
		variable sub_data : STD_LOGIC_VECTOR(1 DOWNTO 0); -- 0 - regs 1 - memory
		variable load_adress : STD_LOGIC_VECTOR(3 DOWNTO 0);
		-- check flag
		variable ready : std_logic;
	BEGIN
		IF (rst = '1') THEN
			ready := '0';
			ready_w <= '0';
			data := (OTHERS => '0');
			valid_map := '0';
			ready_map := '1';
		ELSIF (rising_edge(clk)) THEN
			IF valid_map = '1' THEN
				valid_map := '0';
				ready := '0';
			END IF;

			IF ready_map = '1' AND valid_r = '1' and ready = '0' THEN
				ready_map := '0';
				ready := '1';
				data := data_in; --forming write data
				sub_data := sub_data_in;
				load_adress := load_adr_in;
                if sub_data = "01" then
                    adres_memory <= load_adress;
					memory_data <= data;
                    question_memory <= '1';
                elsif sub_data = "10" or sub_data = "00" then
                    adres_registers <= load_adress;
					registers_data <= data;
                    question_registers <= '1';
                end if;
			END IF;

			IF valid_map = '0' and ready = '1' and (memory_data_ready = '1' or registers_data_ready = '1') then
				valid_map := '1';
				ready_map := '1';
			END IF;
			ready_w <= ready_map;
		END IF;
	END PROCESS; -- main
END rtl; -- rtl